//=========================================================================
// Name & Email must be EXACTLY as in Gradescope roster!
// Name:Garvin Ha 
// Email:gha003@ucr.edu
// 
// Assignment name: Lab2-DatapathControlUnits
// Lab section: 021
// TA: Eren, Omar
// 
// I hereby certify that I have not received assistance on this assignment,
// or used code, from ANY outside source other than the instruction team
// (apart from what was provided in the starter file).
//
//=========================================================================

module aluControlUnit (
    input  wire [1:0] alu_op, 
    input  wire [5:0] instruction_5_0, 
    output reg [3:0] alu_out
    );

// ------------------------------
// Insert your solution below
// ------------------------------ 

endmodule
